.title KiCad schematic
.include "/home/astroelectronica/AE/AP8803/AP8803.spice.txt"
.include "/home/astroelectronica/AE/AP8803/B340B.spice.txt"
.include "/home/astroelectronica/AE/AP8803/WE-TPC.lib"
.include "/home/astroelectronica/AE/AP8803/XPE_SPICE.lib"
.include "/home/astroelectronica/AE/AP8803/c2012x7r2a104k125aa_p.mod"
.include "/home/astroelectronica/AE/AP8803/c3216x7r2a104k160aa_p.mod"
.include "/home/astroelectronica/AE/AP8803/c3225x7r1h475k250ab_p.mod"
D4 /LD3 /LD4 XLampXPEred
R2 VCC /SET {RSET}
D3 /LD2 /LD3 XLampXPEred
D5 /LD4 VCC DI_B340B
XU4 /SET /LD4 C3216X7R2A104K160AA_p
XU5 /LD4 /SW TPC_1038_744066680_68u
D1 /SET /LD1 XLampXPEred
D2 /LD1 /LD2 XLampXPEred
V1 /PWM 0 PULSE(0 {VPUL} {DELAY} {TR} {TF} {DUTY} {CYCLE})
R1 /PWM /CTRL {RCTRL}
XU3 VCC 0 C2012X7R2A104K125AA_p
XU1 /SW  0  /CTRL /SET VCC AL8803_SIMETRIX
V2 VCC 0 {VSOURCE}
XU2 VCC 0 C3225X7R1H475K250AB_p
.end
