.title KiCad schematic
.include "/home/astroelectronica/AE/AP8803/AP8803.spice.txt"
.model __D5 D
D2 /LD2 /LD1 LED
D1 /LD1 /SET LED
R2 VCC /SET R
D3 /LD3 /LD2 LED
D4 /LD4 /LD3 LED
D5 /LD4 VCC __D5
C3 /SET /LD4 C
L1 /LD4 /SW L
C2 VCC 0 C
R1 /PWM /CTRL R
V1 /PWM 0 PULSE( ) 
XU1 NC-U1-0 NC-U1-1 NC-U1-2 NC-U1-3 NC-U1-4 AL8803_SIMETRIX
C1 VCC 0 C
V2 VCC 0 DC {VSOURCE} 
.end
